
//����ת�ã��� 16 �� 64λ���ֻ�ת��Ϊ 64 �� 16λ����λ����
module switch(
	
	input [63:0] patial_product_0,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_1,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_2,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_3,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_4,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_5,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_6,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_7,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_8,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_9,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_10,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_11,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_12,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_13,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_14,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_15,    // ����λ��չ��Ĳ��ֻ�
	input [63:0] patial_product_16,    // ����λ��չ��Ĳ��ֻ�
	output wire[16:0] Tree1,
	output wire[16:0] Tree2,
	output wire[16:0] Tree3,
	output wire[16:0] Tree4,
	output wire[16:0] Tree5,
	output wire[16:0] Tree6,
	output wire[16:0] Tree7,
	output wire[16:0] Tree8,
	output wire[16:0] Tree9,
	output wire[16:0] Tree10,
	output wire[16:0] Tree11,
	output wire[16:0] Tree12,
	output wire[16:0] Tree13,
	output wire[16:0] Tree14,
	output wire[16:0] Tree15,
	output wire[16:0] Tree16,
	output wire[16:0] Tree17,
	output wire[16:0] Tree18,
	output wire[16:0] Tree19,
	output wire[16:0] Tree20,
	output wire[16:0] Tree21,
	output wire[16:0] Tree22,
	output wire[16:0] Tree23,
	output wire[16:0] Tree24,
	output wire[16:0] Tree25,
	output wire[16:0] Tree26,
	output wire[16:0] Tree27,
	output wire[16:0] Tree28,
	output wire[16:0] Tree29,
	output wire[16:0] Tree30,
	output wire[16:0] Tree31,
	output wire[16:0] Tree32,
	output wire[16:0] Tree33,
	output wire[16:0] Tree34,
	output wire[16:0] Tree35,
	output wire[16:0] Tree36,
	output wire[16:0] Tree37,
	output wire[16:0] Tree38,
	output wire[16:0] Tree39,
	output wire[16:0] Tree40,
	output wire[16:0] Tree41,
	output wire[16:0] Tree42,
	output wire[16:0] Tree43,
	output wire[16:0] Tree44,
	output wire[16:0] Tree45,
	output wire[16:0] Tree46,
	output wire[16:0] Tree47,
	output wire[16:0] Tree48,
	output wire[16:0] Tree49,
	output wire[16:0] Tree50,
	output wire[16:0] Tree51,
	output wire[16:0] Tree52,
	output wire[16:0] Tree53,
	output wire[16:0] Tree54,
	output wire[16:0] Tree55,
	output wire[16:0] Tree56,
	output wire[16:0] Tree57,
	output wire[16:0] Tree58,
	output wire[16:0] Tree59,
	output wire[16:0] Tree60,
	output wire[16:0] Tree61,
	output wire[16:0] Tree62,
	output wire[16:0] Tree63,
	output wire[16:0] Tree64
);

assign	Tree1	 =	{patial_product_16	[0],	 patial_product_15	[0],	patial_product_14	[0],	patial_product_13	[0],	patial_product_12	[0],	patial_product_11	[0],	patial_product_10	[0],	patial_product_9	[0],	patial_product_8	[0],	patial_product_7	[0],	patial_product_6	[0],	patial_product_5	[0],	patial_product_4	[0],	patial_product_3	[0],	patial_product_2	[0],	patial_product_1	[0],	patial_product_0	[0]};
assign	Tree2	 =	{patial_product_16	[1],	 patial_product_15	[1],	patial_product_14	[1],	patial_product_13	[1],	patial_product_12	[1],	patial_product_11	[1],	patial_product_10	[1],	patial_product_9	[1],	patial_product_8	[1],	patial_product_7	[1],	patial_product_6	[1],	patial_product_5	[1],	patial_product_4	[1],	patial_product_3	[1],	patial_product_2	[1],	patial_product_1	[1],	patial_product_0	[1]};
assign	Tree3	 =	{patial_product_16	[2],	 patial_product_15	[2],	patial_product_14	[2],	patial_product_13	[2],	patial_product_12	[2],	patial_product_11	[2],	patial_product_10	[2],	patial_product_9	[2],	patial_product_8	[2],	patial_product_7	[2],	patial_product_6	[2],	patial_product_5	[2],	patial_product_4	[2],	patial_product_3	[2],	patial_product_2	[2],	patial_product_1	[2],	patial_product_0	[2]};
assign	Tree4	 =	{patial_product_16	[3],	 patial_product_15	[3],	patial_product_14	[3],	patial_product_13	[3],	patial_product_12	[3],	patial_product_11	[3],	patial_product_10	[3],	patial_product_9	[3],	patial_product_8	[3],	patial_product_7	[3],	patial_product_6	[3],	patial_product_5	[3],	patial_product_4	[3],	patial_product_3	[3],	patial_product_2	[3],	patial_product_1	[3],	patial_product_0	[3]};
assign	Tree5	 =	{patial_product_16	[4],	 patial_product_15	[4],	patial_product_14	[4],	patial_product_13	[4],	patial_product_12	[4],	patial_product_11	[4],	patial_product_10	[4],	patial_product_9	[4],	patial_product_8	[4],	patial_product_7	[4],	patial_product_6	[4],	patial_product_5	[4],	patial_product_4	[4],	patial_product_3	[4],	patial_product_2	[4],	patial_product_1	[4],	patial_product_0	[4]};
assign	Tree6	 =	{patial_product_16	[5],	 patial_product_15	[5],	patial_product_14	[5],	patial_product_13	[5],	patial_product_12	[5],	patial_product_11	[5],	patial_product_10	[5],	patial_product_9	[5],	patial_product_8	[5],	patial_product_7	[5],	patial_product_6	[5],	patial_product_5	[5],	patial_product_4	[5],	patial_product_3	[5],	patial_product_2	[5],	patial_product_1	[5],	patial_product_0	[5]};
assign	Tree7	 =	{patial_product_16	[6],	 patial_product_15	[6],	patial_product_14	[6],	patial_product_13	[6],	patial_product_12	[6],	patial_product_11	[6],	patial_product_10	[6],	patial_product_9	[6],	patial_product_8	[6],	patial_product_7	[6],	patial_product_6	[6],	patial_product_5	[6],	patial_product_4	[6],	patial_product_3	[6],	patial_product_2	[6],	patial_product_1	[6],	patial_product_0	[6]};
assign	Tree8	 =	{patial_product_16	[7],	 patial_product_15	[7],	patial_product_14	[7],	patial_product_13	[7],	patial_product_12	[7],	patial_product_11	[7],	patial_product_10	[7],	patial_product_9	[7],	patial_product_8	[7],	patial_product_7	[7],	patial_product_6	[7],	patial_product_5	[7],	patial_product_4	[7],	patial_product_3	[7],	patial_product_2	[7],	patial_product_1	[7],	patial_product_0	[7]};
assign	Tree9	 =	{patial_product_16	[8],	 patial_product_15	[8],	patial_product_14	[8],	patial_product_13	[8],	patial_product_12	[8],	patial_product_11	[8],	patial_product_10	[8],	patial_product_9	[8],	patial_product_8	[8],	patial_product_7	[8],	patial_product_6	[8],	patial_product_5	[8],	patial_product_4	[8],	patial_product_3	[8],	patial_product_2	[8],	patial_product_1	[8],	patial_product_0	[8]};
assign	Tree10	 =	{patial_product_16	[9],	 patial_product_15	[9],	patial_product_14	[9],	patial_product_13	[9],	patial_product_12	[9],	patial_product_11	[9],	patial_product_10	[9],	patial_product_9	[9],	patial_product_8	[9],	patial_product_7	[9],	patial_product_6	[9],	patial_product_5	[9],	patial_product_4	[9],	patial_product_3	[9],	patial_product_2	[9],	patial_product_1	[9],	patial_product_0	[9]};
assign	Tree11	 =	{patial_product_16	[10],	 patial_product_15	[10],	patial_product_14	[10],	patial_product_13	[10],	patial_product_12	[10],	patial_product_11	[10],	patial_product_10	[10],	patial_product_9	[10],	patial_product_8	[10],	patial_product_7	[10],	patial_product_6	[10],	patial_product_5	[10],	patial_product_4	[10],	patial_product_3	[10],	patial_product_2	[10],	patial_product_1	[10],	patial_product_0	[10]};
assign	Tree12	 =	{patial_product_16	[11],	 patial_product_15	[11],	patial_product_14	[11],	patial_product_13	[11],	patial_product_12	[11],	patial_product_11	[11],	patial_product_10	[11],	patial_product_9	[11],	patial_product_8	[11],	patial_product_7	[11],	patial_product_6	[11],	patial_product_5	[11],	patial_product_4	[11],	patial_product_3	[11],	patial_product_2	[11],	patial_product_1	[11],	patial_product_0	[11]};
assign	Tree13	 =	{patial_product_16	[12],	 patial_product_15	[12],	patial_product_14	[12],	patial_product_13	[12],	patial_product_12	[12],	patial_product_11	[12],	patial_product_10	[12],	patial_product_9	[12],	patial_product_8	[12],	patial_product_7	[12],	patial_product_6	[12],	patial_product_5	[12],	patial_product_4	[12],	patial_product_3	[12],	patial_product_2	[12],	patial_product_1	[12],	patial_product_0	[12]};
assign	Tree14	 =	{patial_product_16	[13],	 patial_product_15	[13],	patial_product_14	[13],	patial_product_13	[13],	patial_product_12	[13],	patial_product_11	[13],	patial_product_10	[13],	patial_product_9	[13],	patial_product_8	[13],	patial_product_7	[13],	patial_product_6	[13],	patial_product_5	[13],	patial_product_4	[13],	patial_product_3	[13],	patial_product_2	[13],	patial_product_1	[13],	patial_product_0	[13]};
assign	Tree15	 =	{patial_product_16	[14],	 patial_product_15	[14],	patial_product_14	[14],	patial_product_13	[14],	patial_product_12	[14],	patial_product_11	[14],	patial_product_10	[14],	patial_product_9	[14],	patial_product_8	[14],	patial_product_7	[14],	patial_product_6	[14],	patial_product_5	[14],	patial_product_4	[14],	patial_product_3	[14],	patial_product_2	[14],	patial_product_1	[14],	patial_product_0	[14]};
assign	Tree16	 =	{patial_product_16	[15],	 patial_product_15	[15],	patial_product_14	[15],	patial_product_13	[15],	patial_product_12	[15],	patial_product_11	[15],	patial_product_10	[15],	patial_product_9	[15],	patial_product_8	[15],	patial_product_7	[15],	patial_product_6	[15],	patial_product_5	[15],	patial_product_4	[15],	patial_product_3	[15],	patial_product_2	[15],	patial_product_1	[15],	patial_product_0	[15]};
assign	Tree17	 =	{patial_product_16	[16],	 patial_product_15	[16],	patial_product_14	[16],	patial_product_13	[16],	patial_product_12	[16],	patial_product_11	[16],	patial_product_10	[16],	patial_product_9	[16],	patial_product_8	[16],	patial_product_7	[16],	patial_product_6	[16],	patial_product_5	[16],	patial_product_4	[16],	patial_product_3	[16],	patial_product_2	[16],	patial_product_1	[16],	patial_product_0	[16]};
assign	Tree18	 =	{patial_product_16	[17],	 patial_product_15	[17],	patial_product_14	[17],	patial_product_13	[17],	patial_product_12	[17],	patial_product_11	[17],	patial_product_10	[17],	patial_product_9	[17],	patial_product_8	[17],	patial_product_7	[17],	patial_product_6	[17],	patial_product_5	[17],	patial_product_4	[17],	patial_product_3	[17],	patial_product_2	[17],	patial_product_1	[17],	patial_product_0	[17]};
assign	Tree19	 =	{patial_product_16	[18],	 patial_product_15	[18],	patial_product_14	[18],	patial_product_13	[18],	patial_product_12	[18],	patial_product_11	[18],	patial_product_10	[18],	patial_product_9	[18],	patial_product_8	[18],	patial_product_7	[18],	patial_product_6	[18],	patial_product_5	[18],	patial_product_4	[18],	patial_product_3	[18],	patial_product_2	[18],	patial_product_1	[18],	patial_product_0	[18]};
assign	Tree20	 =	{patial_product_16	[19],	 patial_product_15	[19],	patial_product_14	[19],	patial_product_13	[19],	patial_product_12	[19],	patial_product_11	[19],	patial_product_10	[19],	patial_product_9	[19],	patial_product_8	[19],	patial_product_7	[19],	patial_product_6	[19],	patial_product_5	[19],	patial_product_4	[19],	patial_product_3	[19],	patial_product_2	[19],	patial_product_1	[19],	patial_product_0	[19]};
assign	Tree21	 =	{patial_product_16	[20],	 patial_product_15	[20],	patial_product_14	[20],	patial_product_13	[20],	patial_product_12	[20],	patial_product_11	[20],	patial_product_10	[20],	patial_product_9	[20],	patial_product_8	[20],	patial_product_7	[20],	patial_product_6	[20],	patial_product_5	[20],	patial_product_4	[20],	patial_product_3	[20],	patial_product_2	[20],	patial_product_1	[20],	patial_product_0	[20]};
assign	Tree22	 =	{patial_product_16	[21],	 patial_product_15	[21],	patial_product_14	[21],	patial_product_13	[21],	patial_product_12	[21],	patial_product_11	[21],	patial_product_10	[21],	patial_product_9	[21],	patial_product_8	[21],	patial_product_7	[21],	patial_product_6	[21],	patial_product_5	[21],	patial_product_4	[21],	patial_product_3	[21],	patial_product_2	[21],	patial_product_1	[21],	patial_product_0	[21]};
assign	Tree23	 =	{patial_product_16	[22],	 patial_product_15	[22],	patial_product_14	[22],	patial_product_13	[22],	patial_product_12	[22],	patial_product_11	[22],	patial_product_10	[22],	patial_product_9	[22],	patial_product_8	[22],	patial_product_7	[22],	patial_product_6	[22],	patial_product_5	[22],	patial_product_4	[22],	patial_product_3	[22],	patial_product_2	[22],	patial_product_1	[22],	patial_product_0	[22]};
assign	Tree24	 =	{patial_product_16	[23],	 patial_product_15	[23],	patial_product_14	[23],	patial_product_13	[23],	patial_product_12	[23],	patial_product_11	[23],	patial_product_10	[23],	patial_product_9	[23],	patial_product_8	[23],	patial_product_7	[23],	patial_product_6	[23],	patial_product_5	[23],	patial_product_4	[23],	patial_product_3	[23],	patial_product_2	[23],	patial_product_1	[23],	patial_product_0	[23]};
assign	Tree25	 =	{patial_product_16	[24],	 patial_product_15	[24],	patial_product_14	[24],	patial_product_13	[24],	patial_product_12	[24],	patial_product_11	[24],	patial_product_10	[24],	patial_product_9	[24],	patial_product_8	[24],	patial_product_7	[24],	patial_product_6	[24],	patial_product_5	[24],	patial_product_4	[24],	patial_product_3	[24],	patial_product_2	[24],	patial_product_1	[24],	patial_product_0	[24]};
assign	Tree26	 =	{patial_product_16	[25],	 patial_product_15	[25],	patial_product_14	[25],	patial_product_13	[25],	patial_product_12	[25],	patial_product_11	[25],	patial_product_10	[25],	patial_product_9	[25],	patial_product_8	[25],	patial_product_7	[25],	patial_product_6	[25],	patial_product_5	[25],	patial_product_4	[25],	patial_product_3	[25],	patial_product_2	[25],	patial_product_1	[25],	patial_product_0	[25]};
assign	Tree27	 =	{patial_product_16	[26],	 patial_product_15	[26],	patial_product_14	[26],	patial_product_13	[26],	patial_product_12	[26],	patial_product_11	[26],	patial_product_10	[26],	patial_product_9	[26],	patial_product_8	[26],	patial_product_7	[26],	patial_product_6	[26],	patial_product_5	[26],	patial_product_4	[26],	patial_product_3	[26],	patial_product_2	[26],	patial_product_1	[26],	patial_product_0	[26]};
assign	Tree28	 =	{patial_product_16	[27],	 patial_product_15	[27],	patial_product_14	[27],	patial_product_13	[27],	patial_product_12	[27],	patial_product_11	[27],	patial_product_10	[27],	patial_product_9	[27],	patial_product_8	[27],	patial_product_7	[27],	patial_product_6	[27],	patial_product_5	[27],	patial_product_4	[27],	patial_product_3	[27],	patial_product_2	[27],	patial_product_1	[27],	patial_product_0	[27]};
assign	Tree29	 =	{patial_product_16	[28],	 patial_product_15	[28],	patial_product_14	[28],	patial_product_13	[28],	patial_product_12	[28],	patial_product_11	[28],	patial_product_10	[28],	patial_product_9	[28],	patial_product_8	[28],	patial_product_7	[28],	patial_product_6	[28],	patial_product_5	[28],	patial_product_4	[28],	patial_product_3	[28],	patial_product_2	[28],	patial_product_1	[28],	patial_product_0	[28]};
assign	Tree30	 =	{patial_product_16	[29],	 patial_product_15	[29],	patial_product_14	[29],	patial_product_13	[29],	patial_product_12	[29],	patial_product_11	[29],	patial_product_10	[29],	patial_product_9	[29],	patial_product_8	[29],	patial_product_7	[29],	patial_product_6	[29],	patial_product_5	[29],	patial_product_4	[29],	patial_product_3	[29],	patial_product_2	[29],	patial_product_1	[29],	patial_product_0	[29]};
assign	Tree31	 =	{patial_product_16	[30],	 patial_product_15	[30],	patial_product_14	[30],	patial_product_13	[30],	patial_product_12	[30],	patial_product_11	[30],	patial_product_10	[30],	patial_product_9	[30],	patial_product_8	[30],	patial_product_7	[30],	patial_product_6	[30],	patial_product_5	[30],	patial_product_4	[30],	patial_product_3	[30],	patial_product_2	[30],	patial_product_1	[30],	patial_product_0	[30]};
assign	Tree32	 =	{patial_product_16	[31],	 patial_product_15	[31],	patial_product_14	[31],	patial_product_13	[31],	patial_product_12	[31],	patial_product_11	[31],	patial_product_10	[31],	patial_product_9	[31],	patial_product_8	[31],	patial_product_7	[31],	patial_product_6	[31],	patial_product_5	[31],	patial_product_4	[31],	patial_product_3	[31],	patial_product_2	[31],	patial_product_1	[31],	patial_product_0	[31]};
assign	Tree33	 =	{patial_product_16	[32],	 patial_product_15	[32],	patial_product_14	[32],	patial_product_13	[32],	patial_product_12	[32],	patial_product_11	[32],	patial_product_10	[32],	patial_product_9	[32],	patial_product_8	[32],	patial_product_7	[32],	patial_product_6	[32],	patial_product_5	[32],	patial_product_4	[32],	patial_product_3	[32],	patial_product_2	[32],	patial_product_1	[32],	patial_product_0	[32]};
assign	Tree34	 =	{patial_product_16	[33],	 patial_product_15	[33],	patial_product_14	[33],	patial_product_13	[33],	patial_product_12	[33],	patial_product_11	[33],	patial_product_10	[33],	patial_product_9	[33],	patial_product_8	[33],	patial_product_7	[33],	patial_product_6	[33],	patial_product_5	[33],	patial_product_4	[33],	patial_product_3	[33],	patial_product_2	[33],	patial_product_1	[33],	patial_product_0	[33]};
assign	Tree35	 =	{patial_product_16	[34],	 patial_product_15	[34],	patial_product_14	[34],	patial_product_13	[34],	patial_product_12	[34],	patial_product_11	[34],	patial_product_10	[34],	patial_product_9	[34],	patial_product_8	[34],	patial_product_7	[34],	patial_product_6	[34],	patial_product_5	[34],	patial_product_4	[34],	patial_product_3	[34],	patial_product_2	[34],	patial_product_1	[34],	patial_product_0	[34]};
assign	Tree36	 =	{patial_product_16	[35],	 patial_product_15	[35],	patial_product_14	[35],	patial_product_13	[35],	patial_product_12	[35],	patial_product_11	[35],	patial_product_10	[35],	patial_product_9	[35],	patial_product_8	[35],	patial_product_7	[35],	patial_product_6	[35],	patial_product_5	[35],	patial_product_4	[35],	patial_product_3	[35],	patial_product_2	[35],	patial_product_1	[35],	patial_product_0	[35]};
assign	Tree37	 =	{patial_product_16	[36],	 patial_product_15	[36],	patial_product_14	[36],	patial_product_13	[36],	patial_product_12	[36],	patial_product_11	[36],	patial_product_10	[36],	patial_product_9	[36],	patial_product_8	[36],	patial_product_7	[36],	patial_product_6	[36],	patial_product_5	[36],	patial_product_4	[36],	patial_product_3	[36],	patial_product_2	[36],	patial_product_1	[36],	patial_product_0	[36]};
assign	Tree38	 =	{patial_product_16	[37],	 patial_product_15	[37],	patial_product_14	[37],	patial_product_13	[37],	patial_product_12	[37],	patial_product_11	[37],	patial_product_10	[37],	patial_product_9	[37],	patial_product_8	[37],	patial_product_7	[37],	patial_product_6	[37],	patial_product_5	[37],	patial_product_4	[37],	patial_product_3	[37],	patial_product_2	[37],	patial_product_1	[37],	patial_product_0	[37]};
assign	Tree39	 =	{patial_product_16	[38],	 patial_product_15	[38],	patial_product_14	[38],	patial_product_13	[38],	patial_product_12	[38],	patial_product_11	[38],	patial_product_10	[38],	patial_product_9	[38],	patial_product_8	[38],	patial_product_7	[38],	patial_product_6	[38],	patial_product_5	[38],	patial_product_4	[38],	patial_product_3	[38],	patial_product_2	[38],	patial_product_1	[38],	patial_product_0	[38]};
assign	Tree40	 =	{patial_product_16	[39],	 patial_product_15	[39],	patial_product_14	[39],	patial_product_13	[39],	patial_product_12	[39],	patial_product_11	[39],	patial_product_10	[39],	patial_product_9	[39],	patial_product_8	[39],	patial_product_7	[39],	patial_product_6	[39],	patial_product_5	[39],	patial_product_4	[39],	patial_product_3	[39],	patial_product_2	[39],	patial_product_1	[39],	patial_product_0	[39]};
assign	Tree41	 =	{patial_product_16	[40],	 patial_product_15	[40],	patial_product_14	[40],	patial_product_13	[40],	patial_product_12	[40],	patial_product_11	[40],	patial_product_10	[40],	patial_product_9	[40],	patial_product_8	[40],	patial_product_7	[40],	patial_product_6	[40],	patial_product_5	[40],	patial_product_4	[40],	patial_product_3	[40],	patial_product_2	[40],	patial_product_1	[40],	patial_product_0	[40]};
assign	Tree42	 =	{patial_product_16	[41],	 patial_product_15	[41],	patial_product_14	[41],	patial_product_13	[41],	patial_product_12	[41],	patial_product_11	[41],	patial_product_10	[41],	patial_product_9	[41],	patial_product_8	[41],	patial_product_7	[41],	patial_product_6	[41],	patial_product_5	[41],	patial_product_4	[41],	patial_product_3	[41],	patial_product_2	[41],	patial_product_1	[41],	patial_product_0	[41]};
assign	Tree43	 =	{patial_product_16	[42],	 patial_product_15	[42],	patial_product_14	[42],	patial_product_13	[42],	patial_product_12	[42],	patial_product_11	[42],	patial_product_10	[42],	patial_product_9	[42],	patial_product_8	[42],	patial_product_7	[42],	patial_product_6	[42],	patial_product_5	[42],	patial_product_4	[42],	patial_product_3	[42],	patial_product_2	[42],	patial_product_1	[42],	patial_product_0	[42]};
assign	Tree44	 =	{patial_product_16	[43],	 patial_product_15	[43],	patial_product_14	[43],	patial_product_13	[43],	patial_product_12	[43],	patial_product_11	[43],	patial_product_10	[43],	patial_product_9	[43],	patial_product_8	[43],	patial_product_7	[43],	patial_product_6	[43],	patial_product_5	[43],	patial_product_4	[43],	patial_product_3	[43],	patial_product_2	[43],	patial_product_1	[43],	patial_product_0	[43]};
assign	Tree45	 =	{patial_product_16	[44],	 patial_product_15	[44],	patial_product_14	[44],	patial_product_13	[44],	patial_product_12	[44],	patial_product_11	[44],	patial_product_10	[44],	patial_product_9	[44],	patial_product_8	[44],	patial_product_7	[44],	patial_product_6	[44],	patial_product_5	[44],	patial_product_4	[44],	patial_product_3	[44],	patial_product_2	[44],	patial_product_1	[44],	patial_product_0	[44]};
assign	Tree46	 =	{patial_product_16	[45],	 patial_product_15	[45],	patial_product_14	[45],	patial_product_13	[45],	patial_product_12	[45],	patial_product_11	[45],	patial_product_10	[45],	patial_product_9	[45],	patial_product_8	[45],	patial_product_7	[45],	patial_product_6	[45],	patial_product_5	[45],	patial_product_4	[45],	patial_product_3	[45],	patial_product_2	[45],	patial_product_1	[45],	patial_product_0	[45]};
assign	Tree47	 =	{patial_product_16	[46],	 patial_product_15	[46],	patial_product_14	[46],	patial_product_13	[46],	patial_product_12	[46],	patial_product_11	[46],	patial_product_10	[46],	patial_product_9	[46],	patial_product_8	[46],	patial_product_7	[46],	patial_product_6	[46],	patial_product_5	[46],	patial_product_4	[46],	patial_product_3	[46],	patial_product_2	[46],	patial_product_1	[46],	patial_product_0	[46]};
assign	Tree48	 =	{patial_product_16	[47],	 patial_product_15	[47],	patial_product_14	[47],	patial_product_13	[47],	patial_product_12	[47],	patial_product_11	[47],	patial_product_10	[47],	patial_product_9	[47],	patial_product_8	[47],	patial_product_7	[47],	patial_product_6	[47],	patial_product_5	[47],	patial_product_4	[47],	patial_product_3	[47],	patial_product_2	[47],	patial_product_1	[47],	patial_product_0	[47]};
assign	Tree49	 =	{patial_product_16	[48],	 patial_product_15	[48],	patial_product_14	[48],	patial_product_13	[48],	patial_product_12	[48],	patial_product_11	[48],	patial_product_10	[48],	patial_product_9	[48],	patial_product_8	[48],	patial_product_7	[48],	patial_product_6	[48],	patial_product_5	[48],	patial_product_4	[48],	patial_product_3	[48],	patial_product_2	[48],	patial_product_1	[48],	patial_product_0	[48]};
assign	Tree50	 =	{patial_product_16	[49],	 patial_product_15	[49],	patial_product_14	[49],	patial_product_13	[49],	patial_product_12	[49],	patial_product_11	[49],	patial_product_10	[49],	patial_product_9	[49],	patial_product_8	[49],	patial_product_7	[49],	patial_product_6	[49],	patial_product_5	[49],	patial_product_4	[49],	patial_product_3	[49],	patial_product_2	[49],	patial_product_1	[49],	patial_product_0	[49]};
assign	Tree51	 =	{patial_product_16	[50],	 patial_product_15	[50],	patial_product_14	[50],	patial_product_13	[50],	patial_product_12	[50],	patial_product_11	[50],	patial_product_10	[50],	patial_product_9	[50],	patial_product_8	[50],	patial_product_7	[50],	patial_product_6	[50],	patial_product_5	[50],	patial_product_4	[50],	patial_product_3	[50],	patial_product_2	[50],	patial_product_1	[50],	patial_product_0	[50]};
assign	Tree52	 =	{patial_product_16	[51],	 patial_product_15	[51],	patial_product_14	[51],	patial_product_13	[51],	patial_product_12	[51],	patial_product_11	[51],	patial_product_10	[51],	patial_product_9	[51],	patial_product_8	[51],	patial_product_7	[51],	patial_product_6	[51],	patial_product_5	[51],	patial_product_4	[51],	patial_product_3	[51],	patial_product_2	[51],	patial_product_1	[51],	patial_product_0	[51]};
assign	Tree53	 =	{patial_product_16	[52],	 patial_product_15	[52],	patial_product_14	[52],	patial_product_13	[52],	patial_product_12	[52],	patial_product_11	[52],	patial_product_10	[52],	patial_product_9	[52],	patial_product_8	[52],	patial_product_7	[52],	patial_product_6	[52],	patial_product_5	[52],	patial_product_4	[52],	patial_product_3	[52],	patial_product_2	[52],	patial_product_1	[52],	patial_product_0	[52]};
assign	Tree54	 =	{patial_product_16	[53],	 patial_product_15	[53],	patial_product_14	[53],	patial_product_13	[53],	patial_product_12	[53],	patial_product_11	[53],	patial_product_10	[53],	patial_product_9	[53],	patial_product_8	[53],	patial_product_7	[53],	patial_product_6	[53],	patial_product_5	[53],	patial_product_4	[53],	patial_product_3	[53],	patial_product_2	[53],	patial_product_1	[53],	patial_product_0	[53]};
assign	Tree55	 =	{patial_product_16	[54],	 patial_product_15	[54],	patial_product_14	[54],	patial_product_13	[54],	patial_product_12	[54],	patial_product_11	[54],	patial_product_10	[54],	patial_product_9	[54],	patial_product_8	[54],	patial_product_7	[54],	patial_product_6	[54],	patial_product_5	[54],	patial_product_4	[54],	patial_product_3	[54],	patial_product_2	[54],	patial_product_1	[54],	patial_product_0	[54]};
assign	Tree56	 =	{patial_product_16	[55],	 patial_product_15	[55],	patial_product_14	[55],	patial_product_13	[55],	patial_product_12	[55],	patial_product_11	[55],	patial_product_10	[55],	patial_product_9	[55],	patial_product_8	[55],	patial_product_7	[55],	patial_product_6	[55],	patial_product_5	[55],	patial_product_4	[55],	patial_product_3	[55],	patial_product_2	[55],	patial_product_1	[55],	patial_product_0	[55]};
assign	Tree57	 =	{patial_product_16	[56],	 patial_product_15	[56],	patial_product_14	[56],	patial_product_13	[56],	patial_product_12	[56],	patial_product_11	[56],	patial_product_10	[56],	patial_product_9	[56],	patial_product_8	[56],	patial_product_7	[56],	patial_product_6	[56],	patial_product_5	[56],	patial_product_4	[56],	patial_product_3	[56],	patial_product_2	[56],	patial_product_1	[56],	patial_product_0	[56]};
assign	Tree58	 =	{patial_product_16	[57],	 patial_product_15	[57],	patial_product_14	[57],	patial_product_13	[57],	patial_product_12	[57],	patial_product_11	[57],	patial_product_10	[57],	patial_product_9	[57],	patial_product_8	[57],	patial_product_7	[57],	patial_product_6	[57],	patial_product_5	[57],	patial_product_4	[57],	patial_product_3	[57],	patial_product_2	[57],	patial_product_1	[57],	patial_product_0	[57]};
assign	Tree59	 =	{patial_product_16	[58],	 patial_product_15	[58],	patial_product_14	[58],	patial_product_13	[58],	patial_product_12	[58],	patial_product_11	[58],	patial_product_10	[58],	patial_product_9	[58],	patial_product_8	[58],	patial_product_7	[58],	patial_product_6	[58],	patial_product_5	[58],	patial_product_4	[58],	patial_product_3	[58],	patial_product_2	[58],	patial_product_1	[58],	patial_product_0	[58]};
assign	Tree60	 =	{patial_product_16	[59],	 patial_product_15	[59],	patial_product_14	[59],	patial_product_13	[59],	patial_product_12	[59],	patial_product_11	[59],	patial_product_10	[59],	patial_product_9	[59],	patial_product_8	[59],	patial_product_7	[59],	patial_product_6	[59],	patial_product_5	[59],	patial_product_4	[59],	patial_product_3	[59],	patial_product_2	[59],	patial_product_1	[59],	patial_product_0	[59]};
assign	Tree61	 =	{patial_product_16	[60],	 patial_product_15	[60],	patial_product_14	[60],	patial_product_13	[60],	patial_product_12	[60],	patial_product_11	[60],	patial_product_10	[60],	patial_product_9	[60],	patial_product_8	[60],	patial_product_7	[60],	patial_product_6	[60],	patial_product_5	[60],	patial_product_4	[60],	patial_product_3	[60],	patial_product_2	[60],	patial_product_1	[60],	patial_product_0	[60]};
assign	Tree62	 =	{patial_product_16	[61],	 patial_product_15	[61],	patial_product_14	[61],	patial_product_13	[61],	patial_product_12	[61],	patial_product_11	[61],	patial_product_10	[61],	patial_product_9	[61],	patial_product_8	[61],	patial_product_7	[61],	patial_product_6	[61],	patial_product_5	[61],	patial_product_4	[61],	patial_product_3	[61],	patial_product_2	[61],	patial_product_1	[61],	patial_product_0	[61]};
assign	Tree63	 =	{patial_product_16	[62],	 patial_product_15	[62],	patial_product_14	[62],	patial_product_13	[62],	patial_product_12	[62],	patial_product_11	[62],	patial_product_10	[62],	patial_product_9	[62],	patial_product_8	[62],	patial_product_7	[62],	patial_product_6	[62],	patial_product_5	[62],	patial_product_4	[62],	patial_product_3	[62],	patial_product_2	[62],	patial_product_1	[62],	patial_product_0	[62]};
assign	Tree64	 =	{patial_product_16	[63],	 patial_product_15	[63],	patial_product_14	[63],	patial_product_13	[63],	patial_product_12	[63],	patial_product_11	[63],	patial_product_10	[63],	patial_product_9	[63],	patial_product_8	[63],	patial_product_7	[63],	patial_product_6	[63],	patial_product_5	[63],	patial_product_4	[63],	patial_product_3	[63],	patial_product_2	[63],	patial_product_1	[63],	patial_product_0	[63]};




endmodule





	